library verilog;
use verilog.vl_types.all;
entity datapath_tb is
end datapath_tb;
