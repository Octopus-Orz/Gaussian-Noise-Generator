library verilog;
use verilog.vl_types.all;
entity MUX_tb is
end MUX_tb;
