library verilog;
use verilog.vl_types.all;
entity LZD_tb is
end LZD_tb;
