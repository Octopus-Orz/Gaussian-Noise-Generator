library verilog;
use verilog.vl_types.all;
entity ROM_trans_new_tb is
end ROM_trans_new_tb;
