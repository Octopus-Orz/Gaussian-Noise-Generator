library verilog;
use verilog.vl_types.all;
entity adder1_tb is
end adder1_tb;
