library verilog;
use verilog.vl_types.all;
entity mult_tb is
end mult_tb;
