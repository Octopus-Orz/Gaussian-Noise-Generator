library verilog;
use verilog.vl_types.all;
entity adder2_tb is
end adder2_tb;
