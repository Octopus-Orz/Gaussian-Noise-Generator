library verilog;
use verilog.vl_types.all;
entity rom_tb is
end rom_tb;
