library verilog;
use verilog.vl_types.all;
entity Mask_tb is
end Mask_tb;
